//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.03 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Fri Dec 20 09:22:35 2024

// addr depth: 1024+1=1025
// data width: 16
// sin tableは1024+1個なので、1024個はSRAMに持って、残りの1つは組み合わせ回路で実現している
module Gowin_pROM_w (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;
wire [15:0] _dout;
wire dff_q_0;

assign gw_gnd = 1'b0;

// ad[10] == 1のとき、16'h7fffを返す
// ad[10] == 0のとき、_doutを返す
// クロックの立ち下がりのときにSRAMが動くので、DFFを使って問題ない。
// DFFには伝搬遅延時間がある、つまりalyawsに影響するのは1サイクル後なので、いい感じになる。

DFFE dff_inst_0 (.Q(dff_q_0), .D(ad[10]), .CLK(clk), .CE(ce));

MUX2 mux_inst_0 (.O(dout[0]), .I0(_dout[0]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_1 (.O(dout[1]), .I0(_dout[1]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_2 (.O(dout[2]), .I0(_dout[2]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_3 (.O(dout[3]), .I0(_dout[3]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_4 (.O(dout[4]), .I0(_dout[4]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_5 (.O(dout[5]), .I0(_dout[5]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_6 (.O(dout[6]), .I0(_dout[6]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_7 (.O(dout[7]), .I0(_dout[7]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_8 (.O(dout[8]), .I0(_dout[8]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_9 (.O(dout[9]), .I0(_dout[9]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_10 (.O(dout[10]), .I0(_dout[10]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_11 (.O(dout[11]), .I0(_dout[11]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_12 (.O(dout[12]), .I0(_dout[12]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_13 (.O(dout[13]), .I0(_dout[13]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_14 (.O(dout[14]), .I0(_dout[14]), .I1(1'd1), .S0(dff_q_0));
MUX2 mux_inst_15 (.O(dout[15]), .I0(_dout[15]), .I1(1'd0), .S0(dff_q_0));

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h02F202C0028D025B022901F701C401920160012E00FB00C90097006500320000;
defparam prom_inst_0.INIT_RAM_01 = 256'h061605E305B1057F054D051B04E804B604840452041F03ED03BB038903560324;
defparam prom_inst_0.INIT_RAM_02 = 256'h0938090608D408A20870083E080C07D907A707750743071106DE06AC067A0648;
defparam prom_inst_0.INIT_RAM_03 = 256'h0C5A0C280BF60BC40B920B600B2D0AFB0AC90A970A650A330A0109CF099D096B;
defparam prom_inst_0.INIT_RAM_04 = 256'h0F790F470F150EE40EB20E800E4E0E1C0DEA0DB80D860D540D220CF00CBE0C8C;
defparam prom_inst_0.INIT_RAM_05 = 256'h129612651233120111CF119E116C113A110810D610A410731041100F0FDD0FAB;
defparam prom_inst_0.INIT_RAM_06 = 256'h15B1157F154D151C14EA14B914871455142413F213C1138F135D132B12FA12C8;
defparam prom_inst_0.INIT_RAM_07 = 256'h18C7189618651833180217D1179F176E173C170B16DA16A816771645161415E2;
defparam prom_inst_0.INIT_RAM_08 = 256'h1BDA1BA91B781B471B161AE51AB41A831A511A2019EF19BE198D195B192A18F9;
defparam prom_inst_0.INIT_RAM_09 = 256'h1EE91EB81E881E571E261DF51DC41D931D621D311D011CD01C9F1C6E1C3D1C0C;
defparam prom_inst_0.INIT_RAM_0A = 256'h21F321C3219221622131210120D0209F206F203E200E1FDD1FAC1F7B1F4B1F1A;
defparam prom_inst_0.INIT_RAM_0B = 256'h24F824C8249824672437240723D723A723762346231622E522B5228422542224;
defparam prom_inst_0.INIT_RAM_0C = 256'h27F727C7279727682738270826D826A826782648261825E825B8258825582528;
defparam prom_inst_0.INIT_RAM_0D = 256'h2AF02AC12A912A622A322A0329D329A429742945291528E528B6288628562827;
defparam prom_inst_0.INIT_RAM_0E = 256'h2DE22DB32D842D552D262CF72CC82C992C6A2C3B2C0C2BDC2BAD2B7E2B4F2B1F;
defparam prom_inst_0.INIT_RAM_0F = 256'h30CD309F3070304230132FE52FB62F872F592F2A2EFB2ECC2E9E2E6F2E402E11;
defparam prom_inst_0.INIT_RAM_10 = 256'h33B133833355332732F932CB329D326E3240321231E431B531873159312A30FC;
defparam prom_inst_0.INIT_RAM_11 = 256'h368D365F3632360435D735A9357B354E352034F234C434973469343B340D33DF;
defparam prom_inst_0.INIT_RAM_12 = 256'h39603933390638D938AC387F3852382537F737CA379D37703742371536E836BA;
defparam prom_inst_0.INIT_RAM_13 = 256'h3C2A3BFE3BD23BA53B793B4C3B203AF33AC63A9A3A6D3A403A1339E739BA398D;
defparam prom_inst_0.INIT_RAM_14 = 256'h3EEC3EC03E943E683E3C3E103DE43DB83D8C3D603D343D083CDC3CAF3C833C57;
defparam prom_inst_0.INIT_RAM_15 = 256'h41A34178414D412140F640CB409F40744048401D3FF13FC63F9A3F6F3F433F17;
defparam prom_inst_0.INIT_RAM_16 = 256'h4450442643FB43D143A6437B4351432642FB42D042A5427A424F422441F941CE;
defparam prom_inst_0.INIT_RAM_17 = 256'h46F346C9469F4675464B462145F745CD45A34579454F452444FA44D044A5447B;
defparam prom_inst_0.INIT_RAM_18 = 256'h498B49624939490F48E648BD4893486A4840481747ED47C4479A47704747471D;
defparam prom_inst_0.INIT_RAM_19 = 256'h4C174BEF4BC74B9E4B754B4D4B244AFB4AD34AAA4A814A584A2F4A0649DD49B4;
defparam prom_inst_0.INIT_RAM_1A = 256'h4E984E714E494E214DF94DD14DA94D814D594D314D094CE14CB94C914C684C40;
defparam prom_inst_0.INIT_RAM_1B = 256'h510D50E650BF50985071504A50234FFB4FD44FAD4F854F5E4F374F0F4EE84EC0;
defparam prom_inst_0.INIT_RAM_1C = 256'h5375534F5329530352DC52B6529052695243521C51F551CF51A85181515B5134;
defparam prom_inst_0.INIT_RAM_1D = 256'h55D055AB55865560553B551554F054CA54A4547F54595433540D53E753C1539B;
defparam prom_inst_0.INIT_RAM_1E = 256'h581E57FA57D557B1578C57675743571E56F956D456AF568A56655640561B55F6;
defparam prom_inst_0.INIT_RAM_1F = 256'h5A5F5A3B5A1859F459D059AC598859645940591C58F858D458B0588C58675843;
defparam prom_inst_0.INIT_RAM_20 = 256'h5C915C6F5C4C5C295C065BE35BC05B9D5B7A5B575B345B105AED5AC95AA65A82;
defparam prom_inst_0.INIT_RAM_21 = 256'h5EB65E945E725E505E2E5E0C5DEA5DC85DA55D835D615D3E5D1C5CF95CD75CB4;
defparam prom_inst_0.INIT_RAM_22 = 256'h60CB60AA608960686047602660055FE45FC25FA15F805F5E5F3C5F1B5EF95ED7;
defparam prom_inst_0.INIT_RAM_23 = 256'h62D262B26292627262526232621161F161D161B06190616F614E612E610D60EC;
defparam prom_inst_0.INIT_RAM_24 = 256'h64CA64AB648B646C644D642E640F63EF63D063B06391637163516332631262F2;
defparam prom_inst_0.INIT_RAM_25 = 256'h66B26693667566576639661B65FC65DE65C065A16582656465456526650764E9;
defparam prom_inst_0.INIT_RAM_26 = 256'h688A686D68506832681567F867DA67BD67A06782676467476729670B66ED66D0;
defparam prom_inst_0.INIT_RAM_27 = 256'h6A526A366A1A69FD69E169C569A9698C697069536937691A68FD68E068C468A7;
defparam prom_inst_0.INIT_RAM_28 = 256'h6C096BEE6BD36BB86B9D6B826B666B4B6B306B146AF86ADD6AC16AA56A896A6E;
defparam prom_inst_0.INIT_RAM_29 = 256'h6DB06D966D7C6D626D486D2E6D146CF96CDF6CC46CAA6C8F6C756C5A6C3F6C24;
defparam prom_inst_0.INIT_RAM_2A = 256'h6F466F2D6F146EFB6EE26EC96EB06E976E7D6E646E4A6E316E176DFE6DE46DCA;
defparam prom_inst_0.INIT_RAM_2B = 256'h70CB70B3709B7083706B7053703B7023700B6FF26FDA6FC26FA96F906F786F5F;
defparam prom_inst_0.INIT_RAM_2C = 256'h723F7228721171FA71E371CC71B5719E7187717071587141712A711270FA70E3;
defparam prom_inst_0.INIT_RAM_2D = 256'h73A0738B7375735F734A7334731E730872F272DC72C572AF72997282726C7255;
defparam prom_inst_0.INIT_RAM_2E = 256'h74F074DC74C774B3749E748974757460744B74367421740B73F673E173CB73B6;
defparam prom_inst_0.INIT_RAM_2F = 256'h762E761B760875F475E175CD75B975A67592757E756A75567542752D75197505;
defparam prom_inst_0.INIT_RAM_30 = 256'h775A774877367723771176FE76EC76D976C776B476A1768E767B766876557642;
defparam prom_inst_0.INIT_RAM_31 = 256'h7874786378517840782F781E780C77FB77E977D877C677B477A27790777E776C;
defparam prom_inst_0.INIT_RAM_32 = 256'h797A796A795B794A793A792A791A790A78F978E978D878C878B778A678957885;
defparam prom_inst_0.INIT_RAM_33 = 256'h7A6E7A607A517A427A337A247A157A0679F779E779D879C979B979AA799A798A;
defparam prom_inst_0.INIT_RAM_34 = 256'h7B507B427B347B277B197B0B7AFD7AEF7AE17AD37AC57AB77AA87A9A7A8C7A7D;
defparam prom_inst_0.INIT_RAM_35 = 256'h7C1E7C117C057BF97BEC7BDF7BD37BC67BB97BAC7B9F7B927B857B787B6A7B5D;
defparam prom_inst_0.INIT_RAM_36 = 256'h7CD97CCE7CC27CB77CAC7CA07C957C897C7E7C727C667C5A7C4E7C427C367C2A;
defparam prom_inst_0.INIT_RAM_37 = 256'h7D817D777D6D7D637D587D4E7D447D3A7D2F7D257D1A7D0F7D057CFA7CEF7CE4;
defparam prom_inst_0.INIT_RAM_38 = 256'h7E157E0C7E037DFB7DF27DE97DE07DD67DCD7DC47DBA7DB17DA77D9E7D947D8A;
defparam prom_inst_0.INIT_RAM_39 = 256'h7E967E8E7E877E7F7E787E707E687E607E587E507E487E3F7E377E2F7E267E1E;
defparam prom_inst_0.INIT_RAM_3A = 256'h7F037EFD7EF77EF07EEA7EE37EDD7ED67ECF7EC87EC17EBA7EB37EAC7EA57E9D;
defparam prom_inst_0.INIT_RAM_3B = 256'h7F5D7F587F537F4E7F497F437F3E7F387F337F2D7F277F227F1C7F167F107F0A;
defparam prom_inst_0.INIT_RAM_3C = 256'h7FA37FA07F9C7F987F947F907F8B7F877F837F7E7F7A7F757F717F6C7F677F62;
defparam prom_inst_0.INIT_RAM_3D = 256'h7FD67FD37FD17FCE7FCB7FC87FC57FC27FBF7FBC7FB97FB57FB27FAE7FAB7FA7;
defparam prom_inst_0.INIT_RAM_3E = 256'h7FF57FF47FF27FF17FEF7FED7FEC7FEA7FE87FE67FE47FE27FE07FDD7FDB7FD9;
defparam prom_inst_0.INIT_RAM_3F = 256'h7FFF7FFF7FFF7FFF7FFF7FFF7FFE7FFE7FFD7FFC7FFB7FFA7FF97FF87FF77FF6;

endmodule //Gowin_pROM_w
